
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "rewind_loop_interface.svh"
`include "rewind_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer2_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer2_out_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer2_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer2_out_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.layer2_out_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.layer2_out_blk_n & AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.layer2_out_blk_n & AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.layer2_out_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer3_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer3_out_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer3_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer3_out_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.layer3_out_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.layer3_out_blk_n);
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer5_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer5_out_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer5_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer5_out_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.layer5_out_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.layer5_out_blk_n);
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer6_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer6_out_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer6_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer6_out_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.layer6_out_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.layer6_out_blk_n);
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer8_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer8_out_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer8_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer8_out_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.layer8_out_blk_n);
    assign fifo_intf_5.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.layer8_out_blk_n);
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer9_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer9_out_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer9_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer9_out_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.layer9_out_blk_n);
    assign fifo_intf_6.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.layer9_out_blk_n);
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer11_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer11_out_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer11_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer11_out_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.layer11_out_blk_n);
    assign fifo_intf_7.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.layer11_out_blk_n);
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer12_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer12_out_U.if_empty_n;
    assign fifo_intf_8.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer12_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer12_out_U.if_full_n;
    assign fifo_intf_8.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.layer12_out_blk_n);
    assign fifo_intf_8.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.layer12_out_blk_n);
    assign fifo_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer14_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer14_out_U.if_empty_n;
    assign fifo_intf_9.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer14_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer14_out_U.if_full_n;
    assign fifo_intf_9.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.layer14_out_blk_n);
    assign fifo_intf_9.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.layer14_out_blk_n);
    assign fifo_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer16_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer16_out_U.if_empty_n;
    assign fifo_intf_10.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer16_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer16_out_U.if_full_n;
    assign fifo_intf_10.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.layer16_out_blk_n);
    assign fifo_intf_10.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.layer16_out_blk_n);
    assign fifo_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_process_data.grp_myproject_fu_7481.layer18_out_U.if_read & AESL_inst_process_data.grp_myproject_fu_7481.layer18_out_U.if_empty_n;
    assign fifo_intf_11.wr_en = AESL_inst_process_data.grp_myproject_fu_7481.layer18_out_U.if_write & AESL_inst_process_data.grp_myproject_fu_7481.layer18_out_U.if_full_n;
    assign fifo_intf_11.fifo_rd_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.grp_softmax_stable_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_s_fu_20.layer18_out_blk_n);
    assign fifo_intf_11.fifo_wr_block = ~(AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.layer18_out_blk_n);
    assign fifo_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_process_data.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_process_data.ap_start == 1'b1 && AESL_inst_process_data.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_process_data.ap_done == 1'b1 && AESL_inst_process_data.ap_continue == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end

logic region_1_idle;
logic [31:0] region_1_start_cnt;
logic [31:0] region_1_done_cnt;
assign region_1_idle = (region_1_start_cnt == region_1_done_cnt) && AESL_inst_process_data.grp_myproject_fu_7481.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_start_cnt <= 32'h0;
    else if (AESL_inst_process_data.grp_myproject_fu_7481.ap_start == 1'b1 && AESL_inst_process_data.grp_myproject_fu_7481.ap_ready == 1'b1)
        region_1_start_cnt <= region_1_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_done_cnt <= 32'h0;
    else if (AESL_inst_process_data.grp_myproject_fu_7481.ap_done == 1'b1 && AESL_inst_process_data.grp_myproject_fu_7481.ap_continue == 1'b1)
        region_1_done_cnt <= region_1_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.real_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.layer2_out_blk_n | ~AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.layer2_out_blk_n | ~AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.layer2_out_blk_n;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_1_idle;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.real_start;
    assign process_intf_2.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.layer2_out_blk_n;
    assign process_intf_2.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.layer3_out_blk_n;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_1_idle;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.real_start;
    assign process_intf_3.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.layer3_out_blk_n;
    assign process_intf_3.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config5_U0.layer5_out_blk_n;
    assign process_intf_3.cin_stall = 1'b0;
    assign process_intf_3.cout_stall = 1'b0;
    assign process_intf_3.region_idle = region_1_idle;
    assign process_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.real_start;
    assign process_intf_4.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.layer5_out_blk_n;
    assign process_intf_4.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.layer6_out_blk_n;
    assign process_intf_4.cin_stall = 1'b0;
    assign process_intf_4.cout_stall = 1'b0;
    assign process_intf_4.region_idle = region_1_idle;
    assign process_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.real_start;
    assign process_intf_5.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.layer6_out_blk_n;
    assign process_intf_5.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.layer8_out_blk_n;
    assign process_intf_5.cin_stall = 1'b0;
    assign process_intf_5.cout_stall = 1'b0;
    assign process_intf_5.region_idle = region_1_idle;
    assign process_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;
    df_process_intf process_intf_6(clock,reset);
    assign process_intf_6.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_start;
    assign process_intf_6.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_ready;
    assign process_intf_6.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_done;
    assign process_intf_6.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_continue;
    assign process_intf_6.real_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.real_start;
    assign process_intf_6.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.layer8_out_blk_n;
    assign process_intf_6.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.layer9_out_blk_n;
    assign process_intf_6.cin_stall = 1'b0;
    assign process_intf_6.cout_stall = 1'b0;
    assign process_intf_6.region_idle = region_1_idle;
    assign process_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_6;
    csv_file_dump pstatus_csv_dumper_6;
    df_process_monitor process_monitor_6;
    df_process_intf process_intf_7(clock,reset);
    assign process_intf_7.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_start;
    assign process_intf_7.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_ready;
    assign process_intf_7.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_done;
    assign process_intf_7.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_continue;
    assign process_intf_7.real_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.real_start;
    assign process_intf_7.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.layer9_out_blk_n;
    assign process_intf_7.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.layer11_out_blk_n;
    assign process_intf_7.cin_stall = 1'b0;
    assign process_intf_7.cout_stall = 1'b0;
    assign process_intf_7.region_idle = region_1_idle;
    assign process_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_7;
    csv_file_dump pstatus_csv_dumper_7;
    df_process_monitor process_monitor_7;
    df_process_intf process_intf_8(clock,reset);
    assign process_intf_8.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_start;
    assign process_intf_8.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_ready;
    assign process_intf_8.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_done;
    assign process_intf_8.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_continue;
    assign process_intf_8.real_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.real_start;
    assign process_intf_8.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.layer11_out_blk_n;
    assign process_intf_8.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.layer12_out_blk_n;
    assign process_intf_8.cin_stall = 1'b0;
    assign process_intf_8.cout_stall = 1'b0;
    assign process_intf_8.region_idle = region_1_idle;
    assign process_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_8;
    csv_file_dump pstatus_csv_dumper_8;
    df_process_monitor process_monitor_8;
    df_process_intf process_intf_9(clock,reset);
    assign process_intf_9.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_start;
    assign process_intf_9.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_ready;
    assign process_intf_9.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_done;
    assign process_intf_9.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_continue;
    assign process_intf_9.real_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.real_start;
    assign process_intf_9.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.layer12_out_blk_n;
    assign process_intf_9.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.layer14_out_blk_n;
    assign process_intf_9.cin_stall = 1'b0;
    assign process_intf_9.cout_stall = 1'b0;
    assign process_intf_9.region_idle = region_1_idle;
    assign process_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_9;
    csv_file_dump pstatus_csv_dumper_9;
    df_process_monitor process_monitor_9;
    df_process_intf process_intf_10(clock,reset);
    assign process_intf_10.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_start;
    assign process_intf_10.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_ready;
    assign process_intf_10.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_done;
    assign process_intf_10.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_continue;
    assign process_intf_10.real_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.real_start;
    assign process_intf_10.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.layer14_out_blk_n;
    assign process_intf_10.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.layer16_out_blk_n;
    assign process_intf_10.cin_stall = 1'b0;
    assign process_intf_10.cout_stall = 1'b0;
    assign process_intf_10.region_idle = region_1_idle;
    assign process_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_10;
    csv_file_dump pstatus_csv_dumper_10;
    df_process_monitor process_monitor_10;
    df_process_intf process_intf_11(clock,reset);
    assign process_intf_11.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.ap_start;
    assign process_intf_11.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.ap_ready;
    assign process_intf_11.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.ap_done;
    assign process_intf_11.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.ap_continue;
    assign process_intf_11.real_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.real_start;
    assign process_intf_11.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.layer16_out_blk_n;
    assign process_intf_11.pout_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.layer18_out_blk_n;
    assign process_intf_11.cin_stall = 1'b0;
    assign process_intf_11.cout_stall = 1'b0;
    assign process_intf_11.region_idle = region_1_idle;
    assign process_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_11;
    csv_file_dump pstatus_csv_dumper_11;
    df_process_monitor process_monitor_11;
    df_process_intf process_intf_12(clock,reset);
    assign process_intf_12.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.ap_start;
    assign process_intf_12.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.ap_ready;
    assign process_intf_12.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.ap_done;
    assign process_intf_12.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.ap_continue;
    assign process_intf_12.real_start = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.ap_start;
    assign process_intf_12.pin_stall = 1'b0 | ~AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.grp_softmax_stable_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_s_fu_20.layer18_out_blk_n;
    assign process_intf_12.pout_stall = 1'b0;
    assign process_intf_12.cin_stall = 1'b0;
    assign process_intf_12.cout_stall = 1'b0;
    assign process_intf_12.region_idle = region_1_idle;
    assign process_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_12;
    csv_file_dump pstatus_csv_dumper_12;
    df_process_monitor process_monitor_12;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_process_data.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_process_data.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_process_data.ap_done;
    assign module_intf_1.ap_continue = AESL_inst_process_data.ap_continue;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.ap_done;
    assign module_intf_9.ap_continue = AESL_inst_process_data.grp_myproject_fu_7481.ap_continue;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_1u_config3_s_fu_95.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_1u_config3_s_fu_95.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_1u_config3_s_fu_95.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_32u_config6_s_fu_1021.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_32u_config6_s_fu_1021.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_32u_config6_s_fu_1021.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1983.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1983.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1983.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_64u_config12_s_fu_1983.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_64u_config12_s_fu_1983.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.call_ln286_shift_line_buffer_array_ap_fixed_16_6_5_3_0_64u_config12_s_fu_1983.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.grp_softmax_stable_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_s_fu_20.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.grp_softmax_stable_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_s_fu_20.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_process_data.grp_myproject_fu_7481.softmax_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_U0.grp_softmax_stable_array_array_ap_fixed_16_6_5_3_0_3u_softmax_config19_s_fu_20.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;

    rewind_loop_intf#(2) rewind_loop_intf_1(clock,reset);
    assign rewind_loop_intf_1.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_1.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_1.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_1.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_enable_reg_pp0_iter0;
    assign rewind_loop_intf_1.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_1.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_1.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_1.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_1.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_1.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_CS_fsm;
    assign rewind_loop_intf_1.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_start;
    assign rewind_loop_intf_1.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_ready;
    assign rewind_loop_intf_1.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config3_s_fu_80.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config3_mult_s_fu_123.ap_done;
    assign rewind_loop_intf_1.loop_continue = 1'b1;
    assign rewind_loop_intf_1.quit_at_end = 1'b1;
    assign rewind_loop_intf_1.finish = finish;
    csv_file_dump rewind_loop_csv_dumper_1;
    rewind_loop_monitor #(2) rewind_loop_monitor_1;
    rewind_loop_intf#(2) rewind_loop_intf_2(clock,reset);
    assign rewind_loop_intf_2.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_2.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_2.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_2.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_enable_reg_pp0_iter0;
    assign rewind_loop_intf_2.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_2.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_2.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_2.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_2.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_2.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_CS_fsm;
    assign rewind_loop_intf_2.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_start;
    assign rewind_loop_intf_2.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_ready;
    assign rewind_loop_intf_2.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config6_s_fu_886.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_mult_s_fu_1793.ap_done;
    assign rewind_loop_intf_2.loop_continue = 1'b1;
    assign rewind_loop_intf_2.quit_at_end = 1'b1;
    assign rewind_loop_intf_2.finish = finish;
    csv_file_dump rewind_loop_csv_dumper_2;
    rewind_loop_monitor #(2) rewind_loop_monitor_2;
    rewind_loop_intf#(2) rewind_loop_intf_3(clock,reset);
    assign rewind_loop_intf_3.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_3.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_3.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_3.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_enable_reg_pp0_iter0;
    assign rewind_loop_intf_3.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_3.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_3.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_3.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_3.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_3.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_CS_fsm;
    assign rewind_loop_intf_3.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_start;
    assign rewind_loop_intf_3.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_ready;
    assign rewind_loop_intf_3.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_64u_config9_s_fu_1718.grp_dense_resource_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config9_mult_s_fu_3523.ap_done;
    assign rewind_loop_intf_3.loop_continue = 1'b1;
    assign rewind_loop_intf_3.quit_at_end = 1'b1;
    assign rewind_loop_intf_3.finish = finish;
    csv_file_dump rewind_loop_csv_dumper_3;
    rewind_loop_monitor #(2) rewind_loop_monitor_3;
    rewind_loop_intf#(2) rewind_loop_intf_4(clock,reset);
    assign rewind_loop_intf_4.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_4.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_4.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_4.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_enable_reg_pp0_iter0;
    assign rewind_loop_intf_4.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_4.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_4.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_4.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_4.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_4.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_CS_fsm;
    assign rewind_loop_intf_4.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_start;
    assign rewind_loop_intf_4.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_ready;
    assign rewind_loop_intf_4.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_16_6_5_3_0_32u_config12_s_fu_1718.grp_dense_resource_ap_fixed_ap_fixed_16_6_5_3_0_config12_mult_s_fu_3523.ap_done;
    assign rewind_loop_intf_4.loop_continue = 1'b1;
    assign rewind_loop_intf_4.quit_at_end = 1'b1;
    assign rewind_loop_intf_4.finish = finish;
    csv_file_dump rewind_loop_csv_dumper_4;
    rewind_loop_monitor #(2) rewind_loop_monitor_4;
    rewind_loop_intf#(2) rewind_loop_intf_5(clock,reset);
    assign rewind_loop_intf_5.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_5.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_5.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_5.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_enable_reg_pp0_iter0;
    assign rewind_loop_intf_5.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_5.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_5.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_5.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_5.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_5.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_CS_fsm;
    assign rewind_loop_intf_5.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_start;
    assign rewind_loop_intf_5.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_ready;
    assign rewind_loop_intf_5.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config16_s_fu_3817.ap_done;
    assign rewind_loop_intf_5.loop_continue = 1'b1;
    assign rewind_loop_intf_5.quit_at_end = 1'b1;
    assign rewind_loop_intf_5.finish = finish;
    csv_file_dump rewind_loop_csv_dumper_5;
    rewind_loop_monitor #(2) rewind_loop_monitor_5;
    rewind_loop_intf#(2) rewind_loop_intf_6(clock,reset);
    assign rewind_loop_intf_6.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_6.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_6.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_ST_fsm_pp0_stage0;
    assign rewind_loop_intf_6.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_enable_reg_pp0_iter0;
    assign rewind_loop_intf_6.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_6.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_6.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_6.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_enable_reg_pp0_iter1;
    assign rewind_loop_intf_6.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_block_pp0_stage0_subdone;
    assign rewind_loop_intf_6.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_CS_fsm;
    assign rewind_loop_intf_6.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_start;
    assign rewind_loop_intf_6.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_ready;
    assign rewind_loop_intf_6.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_8u_array_ap_fixed_16_6_5_3_0_3u_config18_U0.grp_dense_wrapper_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config18_s_fu_67.ap_done;
    assign rewind_loop_intf_6.loop_continue = 1'b1;
    assign rewind_loop_intf_6.quit_at_end = 1'b1;
    assign rewind_loop_intf_6.finish = finish;
    csv_file_dump rewind_loop_csv_dumper_6;
    rewind_loop_monitor #(2) rewind_loop_monitor_6;
    seq_loop_intf#(419) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state37;
    assign seq_loop_intf_1.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.pre_loop_state1 = 419'h0;
    assign seq_loop_intf_1.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state114;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state38;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_process_data.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_process_data.ap_ST_fsm_state38;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_process_data.ap_ST_fsm_state113;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(419) seq_loop_monitor_1;
    seq_loop_intf#(419) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state114;
    assign seq_loop_intf_2.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.pre_loop_state1 = 419'h0;
    assign seq_loop_intf_2.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state37;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state116;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_process_data.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_process_data.ap_ST_fsm_state115;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_process_data.ap_ST_fsm_state267;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(419) seq_loop_monitor_2;
    seq_loop_intf#(419) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state36;
    assign seq_loop_intf_3.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.pre_loop_state1 = 419'h0;
    assign seq_loop_intf_3.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state269;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state37;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_process_data.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_process_data.ap_ST_fsm_state37;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_process_data.ap_ST_fsm_state116;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(419) seq_loop_monitor_3;
    seq_loop_intf#(419) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state36;
    assign seq_loop_intf_4.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.pre_loop_state1 = AESL_inst_process_data.ap_ST_fsm_state343;
    assign seq_loop_intf_4.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state1;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_process_data.ap_ST_fsm_state344;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_process_data.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_process_data.ap_ST_fsm_state344;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_process_data.ap_ST_fsm_state419;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(419) seq_loop_monitor_4;
    seq_loop_intf#(3) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_5.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.pre_loop_state1 = 3'h0;
    assign seq_loop_intf_5.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_5.post_states_valid = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_32u_config3_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(3) seq_loop_monitor_5;
    seq_loop_intf#(3) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_6.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.pre_loop_state1 = 3'h0;
    assign seq_loop_intf_6.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_6.post_states_valid = 1'b1;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_64u_config6_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(3) seq_loop_monitor_6;
    seq_loop_intf#(3) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_7.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.pre_loop_state1 = 3'h0;
    assign seq_loop_intf_7.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_7.post_states_valid = 1'b1;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_64u_config9_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(3) seq_loop_monitor_7;
    seq_loop_intf#(3) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_8.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.pre_loop_state1 = 3'h0;
    assign seq_loop_intf_8.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_8.post_states_valid = 1'b1;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_process_data.grp_myproject_fu_7481.conv_2d_cl_array_ap_fixed_64u_array_ap_fixed_16_6_5_3_0_32u_config12_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(3) seq_loop_monitor_8;
    seq_loop_intf#(5) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_9.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_9.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_9.post_states_valid = 1'b1;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_9.quit_states_valid = 1'b1;
    assign seq_loop_intf_9.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_process_data.grp_myproject_fu_7481.dense_array_ap_fixed_32u_array_ap_fixed_16_6_5_3_0_8u_config16_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(5) seq_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_1.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_1.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_918_4_VITIS_LOOP_920_5_fu_6580.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_first_chan_loop_first_chan_frame_loop_fu_6587.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_frame_chan_loop_fu_6692.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_169_1_fu_6996.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(221) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ST_fsm_state1;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ST_fsm_state221;
    assign upc_loop_intf_5.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ST_fsm_state221;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ST_fsm_state221_blk;
    assign upc_loop_intf_5.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ST_fsm_state221_blk;
    assign upc_loop_intf_5.iter_start_enable = 1'b1;
    assign upc_loop_intf_5.iter_end_enable = 1'b1;
    assign upc_loop_intf_5.quit_enable = 1'b1;
    assign upc_loop_intf_5.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_4_fu_7006.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(221) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_651_2_fu_7021.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_399_1_fu_7251.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadTop_PadTopWidth_fu_22.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadMain_CopyMain_fu_28.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.zeropad2d_cl_array_ap_fixed_1u_array_ap_fixed_16_6_5_3_0_1u_config2_U0.grp_zeropad2d_cl_array_array_ap_fixed_1u_config2_Pipeline_PadBottom_PadBottomWidth_fu_36.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_11.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_11.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_done;
    assign upc_loop_intf_11.loop_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config8_U0.ap_continue;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_12.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_12.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_done;
    assign upc_loop_intf_12.loop_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_64u_config11_U0.ap_continue;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_13.quit_enable = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_13.loop_start = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_done;
    assign upc_loop_intf_13.loop_continue = AESL_inst_process_data.grp_myproject_fu_7481.pooling2d_cl_array_array_ap_fixed_16_6_5_3_0_32u_config14_U0.ap_continue;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;
    upc_loop_intf#(1) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_14.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_14.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_930_6_fu_13031.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(1) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_15.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_15.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_941_8_VITIS_LOOP_943_9_fu_13039.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_16.quit_enable = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_16.loop_start = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_process_data.grp_process_data_Pipeline_VITIS_LOOP_954_10_fu_13047.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);
    pstall_csv_dumper_6 = new("./stalling6.csv");
    pstatus_csv_dumper_6 = new("./status6.csv");
    process_monitor_6 = new(pstall_csv_dumper_6,process_intf_6,pstatus_csv_dumper_6);
    pstall_csv_dumper_7 = new("./stalling7.csv");
    pstatus_csv_dumper_7 = new("./status7.csv");
    process_monitor_7 = new(pstall_csv_dumper_7,process_intf_7,pstatus_csv_dumper_7);
    pstall_csv_dumper_8 = new("./stalling8.csv");
    pstatus_csv_dumper_8 = new("./status8.csv");
    process_monitor_8 = new(pstall_csv_dumper_8,process_intf_8,pstatus_csv_dumper_8);
    pstall_csv_dumper_9 = new("./stalling9.csv");
    pstatus_csv_dumper_9 = new("./status9.csv");
    process_monitor_9 = new(pstall_csv_dumper_9,process_intf_9,pstatus_csv_dumper_9);
    pstall_csv_dumper_10 = new("./stalling10.csv");
    pstatus_csv_dumper_10 = new("./status10.csv");
    process_monitor_10 = new(pstall_csv_dumper_10,process_intf_10,pstatus_csv_dumper_10);
    pstall_csv_dumper_11 = new("./stalling11.csv");
    pstatus_csv_dumper_11 = new("./status11.csv");
    process_monitor_11 = new(pstall_csv_dumper_11,process_intf_11,pstatus_csv_dumper_11);
    pstall_csv_dumper_12 = new("./stalling12.csv");
    pstatus_csv_dumper_12 = new("./status12.csv");
    process_monitor_12 = new(pstall_csv_dumper_12,process_intf_12,pstatus_csv_dumper_12);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);


    rewind_loop_csv_dumper_1 = new("./rewind_loop_status1.csv");
    rewind_loop_monitor_1 = new(rewind_loop_intf_1,rewind_loop_csv_dumper_1);
    rewind_loop_csv_dumper_2 = new("./rewind_loop_status2.csv");
    rewind_loop_monitor_2 = new(rewind_loop_intf_2,rewind_loop_csv_dumper_2);
    rewind_loop_csv_dumper_3 = new("./rewind_loop_status3.csv");
    rewind_loop_monitor_3 = new(rewind_loop_intf_3,rewind_loop_csv_dumper_3);
    rewind_loop_csv_dumper_4 = new("./rewind_loop_status4.csv");
    rewind_loop_monitor_4 = new(rewind_loop_intf_4,rewind_loop_csv_dumper_4);
    rewind_loop_csv_dumper_5 = new("./rewind_loop_status5.csv");
    rewind_loop_monitor_5 = new(rewind_loop_intf_5,rewind_loop_csv_dumper_5);
    rewind_loop_csv_dumper_6 = new("./rewind_loop_status6.csv");
    rewind_loop_monitor_6 = new(rewind_loop_intf_6,rewind_loop_csv_dumper_6);

    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(process_monitor_6);
    sample_manager_inst.add_one_monitor(process_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_8);
    sample_manager_inst.add_one_monitor(process_monitor_9);
    sample_manager_inst.add_one_monitor(process_monitor_10);
    sample_manager_inst.add_one_monitor(process_monitor_11);
    sample_manager_inst.add_one_monitor(process_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(rewind_loop_monitor_1);
    sample_manager_inst.add_one_monitor(rewind_loop_monitor_2);
    sample_manager_inst.add_one_monitor(rewind_loop_monitor_3);
    sample_manager_inst.add_one_monitor(rewind_loop_monitor_4);
    sample_manager_inst.add_one_monitor(rewind_loop_monitor_5);
    sample_manager_inst.add_one_monitor(rewind_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
